module outputGain ( input logic ,
                    input logic signed [15:0] outputGainIn,
                    output logic signed [15:0] outputGainOut);

    always_comb begin
        
    end

endmodule